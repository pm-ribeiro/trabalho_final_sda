library verilog;
use verilog.vl_types.all;
entity final_project_vlg_vec_tst is
end final_project_vlg_vec_tst;
