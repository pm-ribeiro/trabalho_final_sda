library verilog;
use verilog.vl_types.all;
entity final_project is
    port(
        altera_reserved_tms: in     vl_logic;
        altera_reserved_tck: in     vl_logic;
        altera_reserved_tdi: in     vl_logic;
        altera_reserved_tdo: out    vl_logic;
        clock           : in     vl_logic;
        enable          : in     vl_logic;
        addresstest     : out    vl_logic_vector(10 downto 0);
        data            : in     vl_logic_vector(7 downto 0);
        wren            : in     vl_logic;
        q               : out    vl_logic_vector(7 downto 0);
        q2_test         : out    vl_logic_vector(7 downto 0)
    );
end final_project;
